package commons;
// State machine states
typedef enum logic [1:0] {
    IDLE,
    FIRST,
    SECOND
} state_t;
endpackage